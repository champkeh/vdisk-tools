conectix             '�Rvbox  Mac      @       @   x   ���E�ƛ��F��W�q33                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        conectix             '�Rvbox  Mac      @       @   x   ���E�ƛ��F��W�q33                                                                                                                                                                                                                                                                                                                                                                                                                                            